library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package UART_datatypes_pkg is -- same as .h-file in c
	

		
	
end package;

package body UART_datatypes_pkg is -- is the function definition

	

	
end package body;
